LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
------------------------------------------
ENTITY Contador_4Bits IS 
	PORT(
		RELOJ50MHz:IN  STD_LOGIC;
		Contador  :OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END Contador_4Bits;

ARCHITECTURE CODE OF Contador_4Bits IS 

SIGNAL PULSO   :STD_LOGIC;
SIGNAL CUENTA_S:STD_LOGIC_VECTOR(3 DOWNTO 0):="0000";

COMPONENT Un_Hz IS 
	PORT(
		RELOJ_50MHz:IN  STD_LOGIC;
		SALIDA_1HZ :OUT STD_LOGIC
	);
END COMPONENT Un_Hz;

BEGIN

M0: Un_Hz PORT MAP(
	RELOJ_50MHz => RELOJ50MHz,
	SALIDA_1HZ  => Pulso
);

CONTANDO:PROCESS(RELOJ50MHz,CUENTA_S)BEGIN
	IF RELOJ50MHz'EVENT AND RELOJ50MHz='1' THEN
		IF PULSO'EVENT AND PULSO='1' THEN
			IF CUENTA_S = "1111" THEN
				CUENTA_S <= "0000";
			ELSE
				CUENTA_S <= CUENTA_S + "0001";
			END IF;
		END IF;
	END IF;
END PROCESS CONTANDO;

Contador <= CUENTA_S;

END CODE;