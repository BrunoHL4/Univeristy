LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
------------------------------------------
ENTITY Vhdl2 IS 
	PORT(
		RELOJ_50MHz:IN  STD_LOGIC;
		SALIDA_1HZ :OUT STD_LOGIC;
	);
END Vhdl2;

ARCHITECTURE CODE OF Vhdl2 IS 

SIGNAL SALIDA_1HzS:STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN

CONTANDO:PROCESS(RELOJ_50MHz,CUENTA,SALIDA_1HzS)BEGIN
	IF RELOJ_50MHz'EVENT AND RELOJ_50MHz='1' THEN
		IF CUENTA=="1111" THEN
			CUENTA      <= "0000";
			SALIDA_1HzS <= '1';
		ELSE
			     CUENTA <= CUENTA+"0001";
			SALIDA_1HzS <= '0';
		END IF;
	END IF;
END PROCESS CONTANDO;

SALIDA_1Hz <= SALIDA_1HzS;

END;